module MSP430x2xx(Load_en, Clk, Rst, Flags);

// Inputs
input		Load_en;
input 	Clk;
input		Rst;
// Outputs
output   [3:0] Flags;

// Signals
// Registers
// Behavior

MSP430x2xx_block_diagram MSP430x2xx ( 
.Load_en	(Load_en), 
.Clk		(Clk),
.Rst		(Rst),
.Flags	(Flags));
/*hadd halfadder (
a, 
b, 
cout, 
s
);*/


endmodule
