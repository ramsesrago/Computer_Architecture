module mem_cache(address, data);

input address;
output data;


endmodule
